// ./src/top.v

module top();

endmodule //top
